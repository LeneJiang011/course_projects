----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:32:23 06/10/2016 
-- Design Name: 
-- Module Name:    substract - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity substract is
port(
     A:in STD_LOGIC;
	  B:in STD_LOGIC;
	  Cin:in STD_LOGIC;
	  Cout:out STD_LOGIC;
	  s:out STD_LOGIC
	  );
end substract;

architecture Behavioral of substract is

begin
     s<= A XOR (B XOR '1') XOR Cin;
	  Cout<=(Cin AND (A XOR (B XOR '1'))) OR (A AND (B XOR '1'));

end Behavioral;

