----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:11:57 06/17/2016 
-- Design Name: 
-- Module Name:    appa_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity appa_1 is
port(
     a: IN STD_LOGIC;
	  b: IN STD_LOGIC;
	  s: OUT STD_LOGIC
     );

end appa_1;

architecture Behavioral of appa_1 is

begin
     s<=(a OR b);

end Behavioral;

